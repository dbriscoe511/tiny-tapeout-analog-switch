magic
tech sky130A
magscale 1 2
timestamp 1761172680
<< nwell >>
rect -1758 -1897 1758 1897
<< mvpmos >>
rect -1500 -1600 1500 1600
<< mvpdiff >>
rect -1558 1588 -1500 1600
rect -1558 -1588 -1546 1588
rect -1512 -1588 -1500 1588
rect -1558 -1600 -1500 -1588
rect 1500 1588 1558 1600
rect 1500 -1588 1512 1588
rect 1546 -1588 1558 1588
rect 1500 -1600 1558 -1588
<< mvpdiffc >>
rect -1546 -1588 -1512 1588
rect 1512 -1588 1546 1588
<< mvnsubdiff >>
rect -1692 1819 1692 1831
rect -1692 1785 -1584 1819
rect 1584 1785 1692 1819
rect -1692 1773 1692 1785
rect -1692 1723 -1634 1773
rect -1692 -1723 -1680 1723
rect -1646 -1723 -1634 1723
rect 1634 1723 1692 1773
rect -1692 -1773 -1634 -1723
rect 1634 -1723 1646 1723
rect 1680 -1723 1692 1723
rect 1634 -1773 1692 -1723
rect -1692 -1785 1692 -1773
rect -1692 -1819 -1584 -1785
rect 1584 -1819 1692 -1785
rect -1692 -1831 1692 -1819
<< mvnsubdiffcont >>
rect -1584 1785 1584 1819
rect -1680 -1723 -1646 1723
rect 1646 -1723 1680 1723
rect -1584 -1819 1584 -1785
<< poly >>
rect -1500 1681 1500 1697
rect -1500 1647 -1484 1681
rect 1484 1647 1500 1681
rect -1500 1600 1500 1647
rect -1500 -1647 1500 -1600
rect -1500 -1681 -1484 -1647
rect 1484 -1681 1500 -1647
rect -1500 -1697 1500 -1681
<< polycont >>
rect -1484 1647 1484 1681
rect -1484 -1681 1484 -1647
<< locali >>
rect -1680 1785 -1584 1819
rect 1584 1785 1680 1819
rect -1680 1723 -1646 1785
rect 1646 1723 1680 1785
rect -1500 1647 -1484 1681
rect 1484 1647 1500 1681
rect -1546 1588 -1512 1604
rect -1546 -1604 -1512 -1588
rect 1512 1588 1546 1604
rect 1512 -1604 1546 -1588
rect -1500 -1681 -1484 -1647
rect 1484 -1681 1500 -1647
rect -1680 -1785 -1646 -1723
rect 1646 -1785 1680 -1723
rect -1680 -1819 -1584 -1785
rect 1584 -1819 1680 -1785
<< viali >>
rect -1484 1647 1484 1681
rect -1546 -1588 -1512 1588
rect 1512 -1588 1546 1588
rect -1484 -1681 1484 -1647
<< metal1 >>
rect -1496 1681 1496 1687
rect -1496 1647 -1484 1681
rect 1484 1647 1496 1681
rect -1496 1641 1496 1647
rect -1552 1588 -1506 1600
rect -1552 -1588 -1546 1588
rect -1512 -1588 -1506 1588
rect -1552 -1600 -1506 -1588
rect 1506 1588 1552 1600
rect 1506 -1588 1512 1588
rect 1546 -1588 1552 1588
rect 1506 -1600 1552 -1588
rect -1496 -1647 1496 -1641
rect -1496 -1681 -1484 -1647
rect 1484 -1681 1496 -1647
rect -1496 -1687 1496 -1681
<< properties >>
string FIXED_BBOX -1663 -1802 1663 1802
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 16.0 l 15.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
