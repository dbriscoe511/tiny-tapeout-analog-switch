magic
tech sky130A
magscale 1 2
timestamp 1761330451
<< error_s >>
rect 4180 -3020 4190 774
rect 3160 -7980 3166 -7940
<< viali >>
rect 480 -2500 540 140
rect 3820 -2500 3880 140
rect 460 -6520 520 -3880
rect 3780 -6540 3840 -3900
rect 2120 -7960 2380 -7920
rect 3160 -7980 3400 -7940
rect 4740 -7960 5000 -7920
rect 2100 -9800 2360 -9760
rect 3100 -9800 3360 -9760
rect 4700 -9800 4960 -9760
<< metal1 >>
rect 600 720 3800 800
rect 600 560 1640 720
rect 2000 560 3800 720
rect 600 400 3800 560
rect 4400 740 7800 800
rect 4400 580 6580 740
rect 6940 580 7800 740
rect 4400 400 7800 580
rect -600 140 4600 200
rect -600 -2500 480 140
rect 540 -2500 3820 140
rect 3880 -2500 4600 140
rect -600 -2600 4600 -2500
rect 7200 -2600 9200 200
rect -600 -3800 200 -2600
rect 800 -2920 3400 -2800
rect 800 -3340 1620 -2920
rect 2040 -3340 3400 -2920
rect 800 -3600 3400 -3340
rect 4800 -3040 7200 -2800
rect 4800 -3280 6620 -3040
rect 6900 -3280 7200 -3040
rect 4800 -3600 7200 -3280
rect 8400 -3800 9200 -2600
rect -600 -3880 4600 -3800
rect -600 -6520 460 -3880
rect 520 -3900 4600 -3880
rect 520 -6520 3780 -3900
rect -600 -6540 3780 -6520
rect 3840 -6540 4600 -3900
rect -600 -6600 4600 -6540
rect 7200 -6600 9200 -3800
rect 600 -6980 3800 -6800
rect 600 -7140 1640 -6980
rect 2000 -7140 3800 -6980
rect 600 -7200 3800 -7140
rect 4400 -6900 7600 -6800
rect 4400 -7060 6620 -6900
rect 6980 -7060 7600 -6900
rect 4400 -7200 7600 -7060
rect 800 -7440 5060 -7400
rect 800 -7800 5400 -7440
rect 1840 -7920 5200 -7800
rect 1840 -7960 2120 -7920
rect 2380 -7940 4740 -7920
rect 2380 -7960 3080 -7940
rect 1840 -8000 3080 -7960
rect 3400 -7960 4740 -7940
rect 5000 -7960 5200 -7920
rect 3400 -7980 5200 -7960
rect 3160 -8000 5200 -7980
rect 1840 -8140 2080 -8000
rect 1840 -8540 2200 -8140
rect 2240 -8600 2280 -8060
rect 2840 -8140 3080 -8000
rect 2840 -8180 3180 -8140
rect 2310 -8410 2730 -8310
rect 1380 -8840 1580 -8780
rect 2160 -8840 2320 -8600
rect 1380 -8940 2320 -8840
rect 1380 -8980 1580 -8940
rect 2160 -9160 2320 -8940
rect 2630 -8820 2730 -8410
rect 2840 -8540 3200 -8180
rect 3240 -8600 3280 -8080
rect 4340 -8160 4620 -8000
rect 3320 -8560 4200 -8160
rect 4340 -8540 4800 -8160
rect 3180 -8820 3340 -8600
rect 2630 -8920 3340 -8820
rect 1780 -9600 2160 -9200
rect 1780 -9740 2100 -9600
rect 2210 -9650 2240 -9160
rect 2630 -9350 2730 -8920
rect 3180 -9160 3340 -8920
rect 3780 -8790 4200 -8560
rect 4840 -8600 4880 -8060
rect 4920 -8310 5600 -8140
rect 4920 -8540 5180 -8310
rect 2280 -9450 2730 -9350
rect 2900 -9580 3160 -9200
rect 2900 -9740 3080 -9580
rect 3200 -9660 3240 -9160
rect 3280 -9210 3780 -9200
rect 4780 -8820 4940 -8600
rect 5174 -8730 5180 -8540
rect 5600 -8730 5606 -8310
rect 4200 -8940 4940 -8820
rect 4780 -9160 4940 -8940
rect 3280 -9580 4200 -9210
rect 4481 -9580 4762 -9201
rect 4480 -9610 4762 -9580
rect 4480 -9740 4640 -9610
rect 4809 -9640 4847 -9160
rect 5180 -9200 5600 -8730
rect 4900 -9560 5600 -9200
rect 4800 -9647 4847 -9640
rect 4800 -9660 4840 -9647
rect 1780 -9760 5020 -9740
rect 1780 -9800 2100 -9760
rect 2360 -9800 3100 -9760
rect 3360 -9800 4700 -9760
rect 4960 -9800 5020 -9760
rect 1780 -9900 5020 -9800
rect 800 -10300 5400 -9900
<< via1 >>
rect 1640 560 2000 720
rect 6580 580 6940 740
rect 1620 -3340 2040 -2920
rect 6620 -3280 6900 -3040
rect 1640 -7140 2000 -6980
rect 6620 -7060 6980 -6900
rect 3780 -9210 4200 -8790
rect 5180 -8730 5600 -8310
<< metal2 >>
rect 1600 720 2034 747
rect 1600 560 1640 720
rect 2000 560 2034 720
rect 1600 -2920 2034 560
rect 6553 740 6987 797
rect 6553 580 6580 740
rect 6940 580 6987 740
rect 1600 -3340 1620 -2920
rect 2040 -3340 2080 -2920
rect 1600 -3360 2080 -3340
rect 6553 -3040 6987 580
rect 6553 -3280 6620 -3040
rect 6900 -3280 6987 -3040
rect 1600 -6980 2034 -3360
rect 1600 -7140 1640 -6980
rect 2000 -7140 2034 -6980
rect 6553 -6483 6987 -3280
rect 6553 -6900 7017 -6483
rect 6553 -7000 6620 -6900
rect 1600 -9643 2034 -7140
rect 6583 -7060 6620 -7000
rect 6980 -7060 7017 -6900
rect 6583 -7180 7017 -7060
rect 3773 -7614 7017 -7180
rect 3773 -8790 4207 -7614
rect 5203 -8304 5637 -8283
rect 5180 -8310 5637 -8304
rect 5600 -8730 5637 -8310
rect 5180 -8736 5637 -8730
rect 3773 -9210 3780 -8790
rect 4200 -9210 4207 -8790
rect 3773 -9217 4207 -9210
rect 5203 -9643 5637 -8736
rect 1600 -10077 5637 -9643
use sky130_fd_pr__nfet_g5v0d10v5_M3AVYS  XM1
timestamp 1761172680
transform 1 0 5908 0 1 -5162
box -1728 -1858 1728 1858
use sky130_fd_pr__nfet_g5v0d10v5_M3AVYS  XM2
timestamp 1761172680
transform 1 0 2148 0 1 -5202
box -1728 -1858 1728 1858
use sky130_fd_pr__pfet_g5v0d10v5_KUGC3C  XM3
timestamp 1761172680
transform 1 0 5938 0 1 -1123
box -1758 -1897 1758 1897
use sky130_fd_pr__pfet_g5v0d10v5_KUGC3C  XM4
timestamp 1761172680
transform 1 0 2178 0 1 -1163
box -1758 -1897 1758 1897
use sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8  XM5
timestamp 1761172680
transform 1 0 4832 0 1 -9394
box -278 -458 278 458
use sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8  XM6
timestamp 1761172680
transform 1 0 3226 0 1 -9394
box -278 -458 278 458
use sky130_fd_pr__pfet_g5v0d10v5_KLD8Y6  XM7
timestamp 1761172680
transform 1 0 3266 0 1 -8359
box -308 -497 308 497
use sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8  XM8
timestamp 1761172680
transform 1 0 2230 0 1 -9394
box -278 -458 278 458
use sky130_fd_pr__pfet_g5v0d10v5_KLD8Y6  XM9
timestamp 1761172680
transform 1 0 4868 0 1 -8349
box -308 -497 308 497
use sky130_fd_pr__pfet_g5v0d10v5_KLD8Y6  XM10
timestamp 1761172680
transform 1 0 2256 0 1 -8349
box -308 -497 308 497
<< labels >>
flabel metal1 800 -7600 1000 -7400 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 9000 -3400 9200 -3200 0 FreeSans 256 0 0 0 SW_PLUS
port 3 nsew
flabel metal1 800 -10200 1000 -10000 0 FreeSans 256 0 0 0 vss
port 1 nsew
flabel metal1 1380 -8980 1580 -8780 0 FreeSans 256 0 0 0 SW_ON
port 2 nsew
flabel metal1 0 -3400 200 -3200 0 FreeSans 256 0 0 0 SW_MINUS
port 4 nsew
flabel metal2 5203 -10077 5637 -8730 0 FreeSans 1600 0 0 0 gate_dummy
flabel metal2 3773 -7614 7017 -7180 0 FreeSans 1600 0 0 0 gate_main
flabel metal1 2630 -8920 3340 -8820 0 FreeSans 1600 0 0 0 n_tog
<< end >>
