** sch_path: /home/ttuser/Desktop/proj/tiny-tapeout-analog-switch/xschem/analog_switch.sch
.subckt analog_switch vdd vss SW_ON SW_PLUS SW_MINUS
*.PININFO vdd:B vss:B SW_ON:I SW_MINUS:B SW_PLUS:B
XM1 SW_PLUS SW_ON_BUF SW_MINUS SW_MINUS sky130_fd_pr__nfet_g5v0d10v5 L=15 W=16 nf=1 m=1
XM3 SW_MINUS nSW_ON SW_PLUS SW_PLUS sky130_fd_pr__pfet_g5v0d10v5 L=15 W=16 nf=1 m=1
XM2 SW_MINUS nSW_ON SW_MINUS SW_MINUS sky130_fd_pr__nfet_g5v0d10v5 L=15 W=16 nf=1 m=1
XM4 SW_MINUS SW_ON_BUF SW_MINUS SW_MINUS sky130_fd_pr__pfet_g5v0d10v5 L=15 W=16 nf=1 m=1
XM6 SW_ON_BUF net1 vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM7 SW_ON_BUF net1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM8 net1 SW_ON vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM10 net1 SW_ON vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM5 nSW_ON SW_ON_BUF vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM9 nSW_ON SW_ON_BUF vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
.ends
.end
