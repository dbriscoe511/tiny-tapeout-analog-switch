magic
tech sky130A
timestamp 1761172680
<< pwell >>
rect -139 -229 139 229
<< mvnmos >>
rect -25 -100 25 100
<< mvndiff >>
rect -54 94 -25 100
rect -54 -94 -48 94
rect -31 -94 -25 94
rect -54 -100 -25 -94
rect 25 94 54 100
rect 25 -94 31 94
rect 48 -94 54 94
rect 25 -100 54 -94
<< mvndiffc >>
rect -48 -94 -31 94
rect 31 -94 48 94
<< mvpsubdiff >>
rect -121 205 121 211
rect -121 188 -67 205
rect 67 188 121 205
rect -121 182 121 188
rect -121 157 -92 182
rect -121 -157 -115 157
rect -98 -157 -92 157
rect 92 157 121 182
rect -121 -182 -92 -157
rect 92 -157 98 157
rect 115 -157 121 157
rect 92 -182 121 -157
rect -121 -188 121 -182
rect -121 -205 -67 -188
rect 67 -205 121 -188
rect -121 -211 121 -205
<< mvpsubdiffcont >>
rect -67 188 67 205
rect -115 -157 -98 157
rect 98 -157 115 157
rect -67 -205 67 -188
<< poly >>
rect -25 136 25 144
rect -25 119 -17 136
rect 17 119 25 136
rect -25 100 25 119
rect -25 -119 25 -100
rect -25 -136 -17 -119
rect 17 -136 25 -119
rect -25 -144 25 -136
<< polycont >>
rect -17 119 17 136
rect -17 -136 17 -119
<< locali >>
rect -115 188 -67 205
rect 67 188 115 205
rect -115 157 -98 188
rect 98 157 115 188
rect -25 119 -17 136
rect 17 119 25 136
rect -48 94 -31 102
rect -48 -102 -31 -94
rect 31 94 48 102
rect 31 -102 48 -94
rect -25 -136 -17 -119
rect 17 -136 25 -119
rect -115 -188 -98 -157
rect 98 -188 115 -157
rect -115 -205 -67 -188
rect 67 -205 115 -188
<< viali >>
rect -17 119 17 136
rect -48 -94 -31 94
rect 31 -94 48 94
rect -17 -136 17 -119
<< metal1 >>
rect -23 136 23 139
rect -23 119 -17 136
rect 17 119 23 136
rect -23 116 23 119
rect -51 94 -28 100
rect -51 -94 -48 94
rect -31 -94 -28 94
rect -51 -100 -28 -94
rect 28 94 51 100
rect 28 -94 31 94
rect 48 -94 51 94
rect 28 -100 51 -94
rect -23 -119 23 -116
rect -23 -136 -17 -119
rect 17 -136 23 -119
rect -23 -139 23 -136
<< properties >>
string FIXED_BBOX -106 -196 106 196
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 2.0 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
